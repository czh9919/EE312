module NOTGATE(
    input wire a_i1
    output wire b_o
    input wire <.>
    output wire <?>
);

assign b_o=~a_i;
assign <?>=~<.>;

endmodule // NOTGATE


module CONTROL
(
	input [6:0] I_CON,
	output [7:0] O_CON
);
always @(*) begin
	case (I_CON)

end
endmodule //CONTROL
`include "vending_machine_def.v"

module vending_machine (

	clk,							// Clock signal
	reset_n,						// Reset signal (active-low)

	i_input_coin,				// coin is inserted.
	i_select_item,				// item is selected.
	i_trigger_return,			// change-return is triggered

	o_available_item,			// Sign of the item availability
	o_output_item,			// Sign of the item withdrawal
	o_return_coin,				// Sign of the coin return
	stopwatch,
	current_total,
	return_temp,
);

	// Ports Declaration
	// Do not modify the module interface
	input clk;
	input reset_n;

	input [`kNumCoins-1:0] i_input_coin;
	input [`kNumItems-1:0] i_select_item;
	input i_trigger_return;

	output reg [`kNumItems-1:0] o_available_item;
	output reg [`kNumItems-1:0] o_output_item;
	output reg [`kNumCoins-1:0] o_return_coin;

	output [3:0] stopwatch;
	output [`kTotalBits-1:0] current_total;
	output [`kTotalBits-1:0] return_temp;
	// Normally, every output is register,
	//   so that it can provide stable value to the outside.

//////////////////////////////////////////////////////////////////////	/

	//we have to return many coins
	reg [`kCoinBits-1:0] returning_coin_0;
	reg [`kCoinBits-1:0] returning_coin_1;
	reg [`kCoinBits-1:0] returning_coin_2;
	reg block_item_0;
	reg block_item_1;
	//check timeout
	reg [3:0] stopwatch;
	//when return triggered
	reg have_to_return;
	reg  [`kTotalBits-1:0] return_temp;
	reg [`kTotalBits-1:0] temp;
////////////////////////////////////////////////////////////////////////

	// Net constant values (prefix kk & CamelCase)
	// Please refer the wikepedia webpate to know the CamelCase practive of writing.
	// http://en.wikipedia.org/wiki/CamelCase
	// Do not modify the values.
	wire [31:0] kkItemPrice [`kNumItems-1:0];	// Price of each item
	wire [31:0] kkCoinValue [`kNumCoins-1:0];	// Value of each coin
	assign kkItemPrice[0] = 400;
	assign kkItemPrice[1] = 500;
	assign kkItemPrice[2] = 1000;
	assign kkItemPrice[3] = 2000;
	assign kkCoinValue[0] = 100;
	assign kkCoinValue[1] = 500;
	assign kkCoinValue[2] = 1000;


	// NOTE: integer will never be used other than special usages.
	// Only used for loop iteration.
	// You may add more integer variables for loop iteration.
	integer i, j, k,l,m,n;

	// Internal states. You may add your own net & reg variables.
	reg [`kTotalBits-1:0] current_total;
	reg [`kItemBits-1:0] num_items [`kNumItems-1:0];
	reg [`kCoinBits-1:0] num_coins [`kNumCoins-1:0];

	// Next internal states. You may add your own net and reg variables.
	reg [`kTotalBits-1:0] current_total_nxt;
	reg [`kItemBits-1:0] num_items_nxt [`kNumItems-1:0];
	reg [`kCoinBits-1:0] num_coins_nxt [`kNumCoins-1:0];

	// Variables. You may add more your own registers.
	reg [`kTotalBits-1:0] input_total, output_total, return_total_0,return_total_1,return_total_2;


	// Combinational logic for the next states
	always @(*) begin
		// TODO: current_total_nxt
		// You don't have to worry about concurrent activations in each input vector (or array).
		case (i_input_coin)
			3'b001:begin
				current_total_nxt=current_total+100;
				num_coins_nxt[0]=num_coins[0]+1;
			end
			3'b010:begin
				current_total_nxt=current_total+500;
				num_coins_nxt[1]=num_coins[1]+1;
			end
			3'b100:begin
				current_total_nxt=current_total+1000;
				num_coins_nxt[2]=num_coins[2]+1;
			end
		endcase
		case (i_select_item)
			3'b001:begin
				current_total_nxt=current_total-400;
				num_items_nxt[0]=num_items[0]+1;
			end
			3'b010:begin
				current_total_nxt=current_total-500;
				num_items_nxt[1]=num_items[1]+1;
			end
			3'b100:begin
				current_total_nxt=current_total-1000;
				num_items_nxt[2]=num_items[2]+1;
			end 
		endcase



		// Calculate the next current_total state. current_total_nxt =

	end


	// Combinational logic for the outputs
	always @(*) begin
	// TODO: o_available_item
		o_available_item=(current_total_nxt>2000)?4'b1111:(
			(current_total>1000)?4'b0111:(
				(current_total>500)?4'b0011:(
					(current_total>400)?4'b0001:4'b0000
				)
			)
		);
		//$display("HELLO1");
		for (i = 0; i<4; i=i+1) begin
			//!o_available_item[i]=(num_items[i]>=10)?0:(10-num_items[i]);	//10 means sold out
			o_output_item[i]=(num_items[i]>=10)?10:num_items[i];			//10 means sold out
		end
		o_return_coin[0]=(num_coins[0]>=returning_coin_0)?returning_coin_0:num_coins[0];
		o_return_coin[1]=(num_coins[1]>=returning_coin_1)?returning_coin_1:num_coins[1];
		o_return_coin[2]=(num_coins[2]>=returning_coin_2)?returning_coin_2:num_coins[2];
		// TODO: o_output_item
		

	end

	// Sequential circuit to reset or update the states
	always @(posedge clk) begin
		if (!reset_n) begin
			// TODO: reset all states.
			for (i = 0; i<3; i=i+1) begin
				current_total=0;
				o_output_item[i]=0;
				num_coins_nxt[i]=0;
				o_return_coin[i]=0;
			end
		end
		else begin
			// TODO: update all states.
			current_total=current_total_nxt;
		    num_coins[0]=num_coins_nxt[0];
			num_coins[1]=num_coins_nxt[1];
			num_coins[2]=num_coins_nxt[2];
			num_items[0]=num_items_nxt[0];
			num_items[1]=num_items_nxt[1];
			num_items[2]=num_items_nxt[2];
			num_items[3]=num_items_nxt[3];
/////////////////////////////////////////////////////////////////////////

			// decreas stopwatch




			//if you have to return some coins then you have to turn on the bit

		while (current_total>=0&&i_trigger_return==1)
			begin
				if (current_total>=1000)
				begin
					returning_coin_2=returning_coin_2+1;
					current_total=current_total-1000;
				end
				if (current_total>=500)
				begin
					returning_coin_2=returning_coin_1+1;
					current_total=current_total-500;

				end
				if (current_total>=100)
				begin
					returning_coin_2=returning_coin_0+1;
					current_total=current_total-100;
				end
			end

		end		   //update all state end
	end	   //always end

endmodule

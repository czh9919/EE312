module CONTROL (
	input [3:0]
);

endmodule //CONTROL
module NOTGATE(
    input wire a_i
    output wire b_o
    input wire <.>
    output wire <?>
);

assign b_o=~a_i;
assign <?>=~<.>;

endmodule // NOTGATE



module NOTGATE(
    input wire a_i
    output wire b_o
    
);



endmodule // NOTGATE



module NOTGATE(
    input wire a_i1
    output wire b_o

);

assign b_o=~a_i;

endmodule // NOTGATE
// module Adventure (
//     input  wire rstn,
//     input  wire [31:0] I2,
//     input  wire [31:0] I4,
//     output reg 
// );

// endmodule //Adventure
module CONTROL (
	
);

endmodule //CONTROL